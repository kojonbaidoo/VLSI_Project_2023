----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 07.04.2023 13:58:01
-- Design Name: 
-- Module Name: four_bit_divider - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity four_bit_divider is
  Port (
  A,B: in std_logic_vector(3 downto 0);
  Q,R: out std_logic_vector(3 downto 0)
  );
end four_bit_divider;

architecture Behavioral of four_bit_divider is
signal A3,A2,A1,A0: std_logic;
signal B3,B2,B1,B0: std_logic;
signal Y3,Y2,Y1,Y0: std_logic;
signal R3,R2,R1,R0: std_logic;

begin
A3 <= A(3);
A2 <= A(2);
A1 <= A(1);
A0 <= A(0);

B3 <= B(3);
B2 <= B(2);
B1 <= B(1);
B0 <= B(0);

Q <= Y3 & Y2 & Y1 & Y0;
R <= R3 & R2 & R1 & R0;

Y3 <= (A3 and not(A2) and not(A1) and not(A0) and not(B3) and not(B2) and not(B1) and B0) or (A3 and not(A2) and not(A1) and A0 and not(B3) and not(B2) and not(B1) and B0) or (A3 and not(A2) and A1 and not(A0) and not(B3) and not(B2) and not(B1) and B0) or (A3 and not(A2) and A1 and A0 and not(B3) and not(B2) and not(B1) and B0) or (A3 and A2 and not(A1) and not(A0) and not(B3) and not(B2) and not(B1) and B0) or (A3 and A2 and not(A1) and A0 and not(B3) and not(B2) and not(B1) and B0) or (A3 and A2 and A1 and not(A0) and not(B3) and not(B2) and not(B1) and B0) or (A3 and A2 and A1 and A0 and not(B3) and not(B2) and not(B1) and B0);
Y2 <= (not(A3) and A2 and not(A1) and not(A0) and not(B3) and not(B2) and not(B1) and B0) or (not(A3) and A2 and not(A1) and A0 and not(B3) and not(B2) and not(B1) and B0) or (not(A3) and A2 and A1 and not(A0) and not(B3) and not(B2) and not(B1) and B0) or (not(A3) and A2 and A1 and A0 and not(B3) and not(B2) and not(B1) and B0) or (A3 and not(A2) and not(A1) and not(A0) and not(B3) and not(B2) and B1 and not(B0)) or (A3 and not(A2) and not(A1) and A0 and not(B3) and not(B2) and B1 and not(B0)) or (A3 and not(A2) and A1 and not(A0) and not(B3) and not(B2) and B1 and not(B0)) or (A3 and not(A2) and A1 and A0 and not(B3) and not(B2) and B1 and not(B0)) or (A3 and A2 and not(A1) and not(A0) and not(B3) and not(B2) and not(B1) and B0) or (A3 and A2 and not(A1) and not(A0) and not(B3) and not(B2) and B1 and not(B0)) or (A3 and A2 and not(A1) and not(A0) and not(B3) and not(B2) and B1 and B0) or (A3 and A2 and not(A1) and A0 and not(B3) and not(B2) and not(B1) and B0) or (A3 and A2 and not(A1) and A0 and not(B3) and not(B2) and B1 and not(B0)) or (A3 and A2 and not(A1) and A0 and not(B3) and not(B2) and B1 and B0) or (A3 and A2 and A1 and not(A0) and not(B3) and not(B2) and not(B1) and B0) or (A3 and A2 and A1 and not(A0) and not(B3) and not(B2) and B1 and not(B0)) or (A3 and A2 and A1 and not(A0) and not(B3) and not(B2) and B1 and B0) or (A3 and A2 and A1 and A0 and not(B3) and not(B2) and not(B1) and B0) or (A3 and A2 and A1 and A0 and not(B3) and not(B2) and B1 and not(B0)) or (A3 and A2 and A1 and A0 and not(B3) and not(B2) and B1 and B0);
Y1 <= (not(A3) and not(A2) and A1 and not(A0) and not(B3) and not(B2) and not(B1) and B0) or (not(A3) and not(A2) and A1 and A0 and not(B3) and not(B2) and not(B1) and B0) or (not(A3) and A2 and not(A1) and not(A0) and not(B3) and not(B2) and B1 and not(B0)) or (not(A3) and A2 and not(A1) and A0 and not(B3) and not(B2) and B1 and not(B0)) or (not(A3) and A2 and A1 and not(A0) and not(B3) and not(B2) and not(B1) and B0) or (not(A3) and A2 and A1 and not(A0) and not(B3) and not(B2) and B1 and not(B0)) or (not(A3) and A2 and A1 and not(A0) and not(B3) and not(B2) and B1 and B0) or (not(A3) and A2 and A1 and A0 and not(B3) and not(B2) and not(B1) and B0) or (not(A3) and A2 and A1 and A0 and not(B3) and not(B2) and B1 and not(B0)) or (not(A3) and A2 and A1 and A0 and not(B3) and not(B2) and B1 and B0) or (A3 and not(A2) and not(A1) and not(A0) and not(B3) and not(B2) and B1 and B0) or (A3 and not(A2) and not(A1) and not(A0) and not(B3) and B2 and not(B1) and not(B0)) or (A3 and not(A2) and not(A1) and A0 and not(B3) and not(B2) and B1 and B0) or (A3 and not(A2) and not(A1) and A0 and not(B3) and B2 and not(B1) and not(B0)) or (A3 and not(A2) and A1 and not(A0) and not(B3) and not(B2) and not(B1) and B0) or (A3 and not(A2) and A1 and not(A0) and not(B3) and not(B2) and B1 and B0) or (A3 and not(A2) and A1 and not(A0) and not(B3) and B2 and not(B1) and not(B0)) or (A3 and not(A2) and A1 and not(A0) and not(B3) and B2 and not(B1) and B0) or (A3 and not(A2) and A1 and A0 and not(B3) and not(B2) and not(B1) and B0) or (A3 and not(A2) and A1 and A0 and not(B3) and not(B2) and B1 and B0) or (A3 and not(A2) and A1 and A0 and not(B3) and B2 and not(B1) and not(B0)) or (A3 and not(A2) and A1 and A0 and not(B3) and B2 and not(B1) and B0) or (A3 and A2 and not(A1) and not(A0) and not(B3) and not(B2) and B1 and not(B0)) or (A3 and A2 and not(A1) and not(A0) and not(B3) and B2 and not(B1) and not(B0)) or (A3 and A2 and not(A1) and not(A0) and not(B3) and B2 and not(B1) and B0) or (A3 and A2 and not(A1) and not(A0) and not(B3) and B2 and B1 and not(B0)) or (A3 and A2 and not(A1) and A0 and not(B3) and not(B2) and B1 and not(B0)) or (A3 and A2 and not(A1) and A0 and not(B3) and B2 and not(B1) and not(B0)) or (A3 and A2 and not(A1) and A0 and not(B3) and B2 and not(B1) and B0) or (A3 and A2 and not(A1) and A0 and not(B3) and B2 and B1 and not(B0)) or (A3 and A2 and A1 and not(A0) and not(B3) and not(B2) and not(B1) and B0) or (A3 and A2 and A1 and not(A0) and not(B3) and not(B2) and B1 and not(B0)) or (A3 and A2 and A1 and not(A0) and not(B3) and B2 and not(B1) and not(B0)) or (A3 and A2 and A1 and not(A0) and not(B3) and B2 and not(B1) and B0) or (A3 and A2 and A1 and not(A0) and not(B3) and B2 and B1 and not(B0)) or (A3 and A2 and A1 and not(A0) and not(B3) and B2 and B1 and B0) or (A3 and A2 and A1 and A0 and not(B3) and not(B2) and not(B1) and B0) or (A3 and A2 and A1 and A0 and not(B3) and not(B2) and B1 and not(B0)) or (A3 and A2 and A1 and A0 and not(B3) and B2 and not(B1) and not(B0)) or (A3 and A2 and A1 and A0 and not(B3) and B2 and not(B1) and B0) or (A3 and A2 and A1 and A0 and not(B3) and B2 and B1 and not(B0)) or (A3 and A2 and A1 and A0 and not(B3) and B2 and B1 and B0);
Y0 <= (not(A3) and not(A2) and not(A1) and A0 and not(B3) and not(B2) and not(B1) and B0) or (not(A3) and not(A2) and A1 and not(A0) and not(B3) and not(B2) and B1 and not(B0)) or (not(A3) and not(A2) and A1 and A0 and not(B3) and not(B2) and not(B1) and B0) or (not(A3) and not(A2) and A1 and A0 and not(B3) and not(B2) and B1 and not(B0)) or (not(A3) and not(A2) and A1 and A0 and not(B3) and not(B2) and B1 and B0) or (not(A3) and A2 and not(A1) and not(A0) and not(B3) and not(B2) and B1 and B0) or (not(A3) and A2 and not(A1) and not(A0) and not(B3) and B2 and not(B1) and not(B0)) or (not(A3) and A2 and not(A1) and A0 and not(B3) and not(B2) and not(B1) and B0) or (not(A3) and A2 and not(A1) and A0 and not(B3) and not(B2) and B1 and B0) or (not(A3) and A2 and not(A1) and A0 and not(B3) and B2 and not(B1) and not(B0)) or (not(A3) and A2 and not(A1) and A0 and not(B3) and B2 and not(B1) and B0) or (not(A3) and A2 and A1 and not(A0) and not(B3) and not(B2) and B1 and not(B0)) or (not(A3) and A2 and A1 and not(A0) and not(B3) and B2 and not(B1) and not(B0)) or (not(A3) and A2 and A1 and not(A0) and not(B3) and B2 and not(B1) and B0) or (not(A3) and A2 and A1 and not(A0) and not(B3) and B2 and B1 and not(B0)) or (not(A3) and A2 and A1 and A0 and not(B3) and not(B2) and not(B1) and B0) or (not(A3) and A2 and A1 and A0 and not(B3) and not(B2) and B1 and not(B0)) or (not(A3) and A2 and A1 and A0 and not(B3) and B2 and not(B1) and not(B0)) or (not(A3) and A2 and A1 and A0 and not(B3) and B2 and not(B1) and B0) or (not(A3) and A2 and A1 and A0 and not(B3) and B2 and B1 and not(B0)) or (not(A3) and A2 and A1 and A0 and not(B3) and B2 and B1 and B0) or (A3 and not(A2) and not(A1) and not(A0) and not(B3) and B2 and not(B1) and B0) or (A3 and not(A2) and not(A1) and not(A0) and not(B3) and B2 and B1 and not(B0)) or (A3 and not(A2) and not(A1) and not(A0) and not(B3) and B2 and B1 and B0) or (A3 and not(A2) and not(A1) and not(A0) and B3 and not(B2) and not(B1) and not(B0)) or (A3 and not(A2) and not(A1) and A0 and not(B3) and not(B2) and not(B1) and B0) or (A3 and not(A2) and not(A1) and A0 and not(B3) and not(B2) and B1 and B0) or (A3 and not(A2) and not(A1) and A0 and not(B3) and B2 and not(B1) and B0) or (A3 and not(A2) and not(A1) and A0 and not(B3) and B2 and B1 and not(B0)) or (A3 and not(A2) and not(A1) and A0 and not(B3) and B2 and B1 and B0) or (A3 and not(A2) and not(A1) and A0 and B3 and not(B2) and not(B1) and not(B0)) or (A3 and not(A2) and not(A1) and A0 and B3 and not(B2) and not(B1) and B0) or (A3 and not(A2) and A1 and not(A0) and not(B3) and not(B2) and B1 and not(B0)) or (A3 and not(A2) and A1 and not(A0) and not(B3) and not(B2) and B1 and B0) or (A3 and not(A2) and A1 and not(A0) and not(B3) and B2 and B1 and not(B0)) or (A3 and not(A2) and A1 and not(A0) and not(B3) and B2 and B1 and B0) or (A3 and not(A2) and A1 and not(A0) and B3 and not(B2) and not(B1) and not(B0)) or (A3 and not(A2) and A1 and not(A0) and B3 and not(B2) and not(B1) and B0) or (A3 and not(A2) and A1 and not(A0) and B3 and not(B2) and B1 and not(B0)) or (A3 and not(A2) and A1 and A0 and not(B3) and not(B2) and not(B1) and B0) or (A3 and not(A2) and A1 and A0 and not(B3) and not(B2) and B1 and not(B0)) or (A3 and not(A2) and A1 and A0 and not(B3) and not(B2) and B1 and B0) or (A3 and not(A2) and A1 and A0 and not(B3) and B2 and B1 and not(B0)) or (A3 and not(A2) and A1 and A0 and not(B3) and B2 and B1 and B0) or (A3 and not(A2) and A1 and A0 and B3 and not(B2) and not(B1) and not(B0)) or (A3 and not(A2) and A1 and A0 and B3 and not(B2) and not(B1) and B0) or (A3 and not(A2) and A1 and A0 and B3 and not(B2) and B1 and not(B0)) or (A3 and not(A2) and A1 and A0 and B3 and not(B2) and B1 and B0) or (A3 and A2 and not(A1) and not(A0) and not(B3) and B2 and not(B1) and not(B0)) or (A3 and A2 and not(A1) and not(A0) and not(B3) and B2 and B1 and B0) or (A3 and A2 and not(A1) and not(A0) and B3 and not(B2) and not(B1) and not(B0)) or (A3 and A2 and not(A1) and not(A0) and B3 and not(B2) and not(B1) and B0) or (A3 and A2 and not(A1) and not(A0) and B3 and not(B2) and B1 and not(B0)) or (A3 and A2 and not(A1) and not(A0) and B3 and not(B2) and B1 and B0) or (A3 and A2 and not(A1) and not(A0) and B3 and B2 and not(B1) and not(B0)) or (A3 and A2 and not(A1) and A0 and not(B3) and not(B2) and not(B1) and B0) or (A3 and A2 and not(A1) and A0 and not(B3) and B2 and not(B1) and not(B0)) or (A3 and A2 and not(A1) and A0 and not(B3) and B2 and B1 and B0) or (A3 and A2 and not(A1) and A0 and B3 and not(B2) and not(B1) and not(B0)) or (A3 and A2 and not(A1) and A0 and B3 and not(B2) and not(B1) and B0) or (A3 and A2 and not(A1) and A0 and B3 and not(B2) and B1 and not(B0)) or (A3 and A2 and not(A1) and A0 and B3 and not(B2) and B1 and B0) or (A3 and A2 and not(A1) and A0 and B3 and B2 and not(B1) and not(B0)) or (A3 and A2 and not(A1) and A0 and B3 and B2 and not(B1) and B0) or (A3 and A2 and A1 and not(A0) and not(B3) and not(B2) and B1 and not(B0)) or (A3 and A2 and A1 and not(A0) and not(B3) and B2 and not(B1) and not(B0)) or (A3 and A2 and A1 and not(A0) and B3 and not(B2) and not(B1) and not(B0)) or (A3 and A2 and A1 and not(A0) and B3 and not(B2) and not(B1) and B0) or (A3 and A2 and A1 and not(A0) and B3 and not(B2) and B1 and not(B0)) or (A3 and A2 and A1 and not(A0) and B3 and not(B2) and B1 and B0) or (A3 and A2 and A1 and not(A0) and B3 and B2 and not(B1) and not(B0)) or (A3 and A2 and A1 and not(A0) and B3 and B2 and not(B1) and B0) or (A3 and A2 and A1 and not(A0) and B3 and B2 and B1 and not(B0)) or (A3 and A2 and A1 and A0 and not(B3) and not(B2) and not(B1) and B0) or (A3 and A2 and A1 and A0 and not(B3) and not(B2) and B1 and not(B0)) or (A3 and A2 and A1 and A0 and not(B3) and not(B2) and B1 and B0) or (A3 and A2 and A1 and A0 and not(B3) and B2 and not(B1) and not(B0)) or (A3 and A2 and A1 and A0 and not(B3) and B2 and not(B1) and B0) or (A3 and A2 and A1 and A0 and B3 and not(B2) and not(B1) and not(B0)) or (A3 and A2 and A1 and A0 and B3 and not(B2) and not(B1) and B0) or (A3 and A2 and A1 and A0 and B3 and not(B2) and B1 and not(B0)) or (A3 and A2 and A1 and A0 and B3 and not(B2) and B1 and B0) or (A3 and A2 and A1 and A0 and B3 and B2 and not(B1) and not(B0)) or (A3 and A2 and A1 and A0 and B3 and B2 and not(B1) and B0) or (A3 and A2 and A1 and A0 and B3 and B2 and B1 and not(B0)) or (A3 and A2 and A1 and A0 and B3 and B2 and B1 and B0);

R3 <= (A3 and not(A2) and not(A1) and not(A0) and B3 and not(B2) and not(B1) and B0) or (A3 and not(A2) and not(A1) and not(A0) and B3 and not(B2) and B1 and not(B0)) or (A3 and not(A2) and not(A1) and not(A0) and B3 and not(B2) and B1 and B0) or (A3 and not(A2) and not(A1) and not(A0) and B3 and B2 and not(B1) and not(B0)) or (A3 and not(A2) and not(A1) and not(A0) and B3 and B2 and not(B1) and B0) or (A3 and not(A2) and not(A1) and not(A0) and B3 and B2 and B1 and not(B0)) or (A3 and not(A2) and not(A1) and not(A0) and B3 and B2 and B1 and B0) or (A3 and not(A2) and not(A1) and A0 and B3 and not(B2) and B1 and not(B0)) or (A3 and not(A2) and not(A1) and A0 and B3 and not(B2) and B1 and B0) or (A3 and not(A2) and not(A1) and A0 and B3 and B2 and not(B1) and not(B0)) or (A3 and not(A2) and not(A1) and A0 and B3 and B2 and not(B1) and B0) or (A3 and not(A2) and not(A1) and A0 and B3 and B2 and B1 and not(B0)) or (A3 and not(A2) and not(A1) and A0 and B3 and B2 and B1 and B0) or (A3 and not(A2) and A1 and not(A0) and B3 and not(B2) and B1 and B0) or (A3 and not(A2) and A1 and not(A0) and B3 and B2 and not(B1) and not(B0)) or (A3 and not(A2) and A1 and not(A0) and B3 and B2 and not(B1) and B0) or (A3 and not(A2) and A1 and not(A0) and B3 and B2 and B1 and not(B0)) or (A3 and not(A2) and A1 and not(A0) and B3 and B2 and B1 and B0) or (A3 and not(A2) and A1 and A0 and B3 and B2 and not(B1) and not(B0)) or (A3 and not(A2) and A1 and A0 and B3 and B2 and not(B1) and B0) or (A3 and not(A2) and A1 and A0 and B3 and B2 and B1 and not(B0)) or (A3 and not(A2) and A1 and A0 and B3 and B2 and B1 and B0) or (A3 and A2 and not(A1) and not(A0) and B3 and B2 and not(B1) and B0) or (A3 and A2 and not(A1) and not(A0) and B3 and B2 and B1 and not(B0)) or (A3 and A2 and not(A1) and not(A0) and B3 and B2 and B1 and B0) or (A3 and A2 and not(A1) and A0 and B3 and B2 and B1 and not(B0)) or (A3 and A2 and not(A1) and A0 and B3 and B2 and B1 and B0) or (A3 and A2 and A1 and not(A0) and B3 and B2 and B1 and B0);
R2 <= (not(A3) and A2 and not(A1) and not(A0) and not(B3) and B2 and not(B1) and B0) or (not(A3) and A2 and not(A1) and not(A0) and not(B3) and B2 and B1 and not(B0)) or (not(A3) and A2 and not(A1) and not(A0) and not(B3) and B2 and B1 and B0) or (not(A3) and A2 and not(A1) and not(A0) and B3 and not(B2) and not(B1) and not(B0)) or (not(A3) and A2 and not(A1) and not(A0) and B3 and not(B2) and not(B1) and B0) or (not(A3) and A2 and not(A1) and not(A0) and B3 and not(B2) and B1 and not(B0)) or (not(A3) and A2 and not(A1) and not(A0) and B3 and not(B2) and B1 and B0) or (not(A3) and A2 and not(A1) and not(A0) and B3 and B2 and not(B1) and not(B0)) or (not(A3) and A2 and not(A1) and not(A0) and B3 and B2 and not(B1) and B0) or (not(A3) and A2 and not(A1) and not(A0) and B3 and B2 and B1 and not(B0)) or (not(A3) and A2 and not(A1) and not(A0) and B3 and B2 and B1 and B0) or (not(A3) and A2 and not(A1) and A0 and not(B3) and B2 and B1 and not(B0)) or (not(A3) and A2 and not(A1) and A0 and not(B3) and B2 and B1 and B0) or (not(A3) and A2 and not(A1) and A0 and B3 and not(B2) and not(B1) and not(B0)) or (not(A3) and A2 and not(A1) and A0 and B3 and not(B2) and not(B1) and B0) or (not(A3) and A2 and not(A1) and A0 and B3 and not(B2) and B1 and not(B0)) or (not(A3) and A2 and not(A1) and A0 and B3 and not(B2) and B1 and B0) or (not(A3) and A2 and not(A1) and A0 and B3 and B2 and not(B1) and not(B0)) or (not(A3) and A2 and not(A1) and A0 and B3 and B2 and not(B1) and B0) or (not(A3) and A2 and not(A1) and A0 and B3 and B2 and B1 and not(B0)) or (not(A3) and A2 and not(A1) and A0 and B3 and B2 and B1 and B0) or (not(A3) and A2 and A1 and not(A0) and not(B3) and B2 and B1 and B0) or (not(A3) and A2 and A1 and not(A0) and B3 and not(B2) and not(B1) and not(B0)) or (not(A3) and A2 and A1 and not(A0) and B3 and not(B2) and not(B1) and B0) or (not(A3) and A2 and A1 and not(A0) and B3 and not(B2) and B1 and not(B0)) or (not(A3) and A2 and A1 and not(A0) and B3 and not(B2) and B1 and B0) or (not(A3) and A2 and A1 and not(A0) and B3 and B2 and not(B1) and not(B0)) or (not(A3) and A2 and A1 and not(A0) and B3 and B2 and not(B1) and B0) or (not(A3) and A2 and A1 and not(A0) and B3 and B2 and B1 and not(B0)) or (not(A3) and A2 and A1 and not(A0) and B3 and B2 and B1 and B0) or (not(A3) and A2 and A1 and A0 and B3 and not(B2) and not(B1) and not(B0)) or (not(A3) and A2 and A1 and A0 and B3 and not(B2) and not(B1) and B0) or (not(A3) and A2 and A1 and A0 and B3 and not(B2) and B1 and not(B0)) or (not(A3) and A2 and A1 and A0 and B3 and not(B2) and B1 and B0) or (not(A3) and A2 and A1 and A0 and B3 and B2 and not(B1) and not(B0)) or (not(A3) and A2 and A1 and A0 and B3 and B2 and not(B1) and B0) or (not(A3) and A2 and A1 and A0 and B3 and B2 and B1 and not(B0)) or (not(A3) and A2 and A1 and A0 and B3 and B2 and B1 and B0) or (A3 and not(A2) and not(A1) and A0 and not(B3) and B2 and not(B1) and B0) or (A3 and not(A2) and A1 and not(A0) and not(B3) and B2 and B1 and not(B0)) or (A3 and not(A2) and A1 and A0 and not(B3) and B2 and B1 and not(B0)) or (A3 and not(A2) and A1 and A0 and not(B3) and B2 and B1 and B0) or (A3 and A2 and not(A1) and not(A0) and not(B3) and B2 and B1 and B0) or (A3 and A2 and not(A1) and not(A0) and B3 and not(B2) and not(B1) and not(B0)) or (A3 and A2 and not(A1) and not(A0) and B3 and B2 and not(B1) and B0) or (A3 and A2 and not(A1) and not(A0) and B3 and B2 and B1 and not(B0)) or (A3 and A2 and not(A1) and not(A0) and B3 and B2 and B1 and B0) or (A3 and A2 and not(A1) and A0 and not(B3) and B2 and B1 and B0) or (A3 and A2 and not(A1) and A0 and B3 and not(B2) and not(B1) and not(B0)) or (A3 and A2 and not(A1) and A0 and B3 and not(B2) and not(B1) and B0) or (A3 and A2 and not(A1) and A0 and B3 and B2 and B1 and not(B0)) or (A3 and A2 and not(A1) and A0 and B3 and B2 and B1 and B0) or (A3 and A2 and A1 and not(A0) and not(B3) and B2 and not(B1) and B0) or (A3 and A2 and A1 and not(A0) and B3 and not(B2) and not(B1) and not(B0)) or (A3 and A2 and A1 and not(A0) and B3 and not(B2) and not(B1) and B0) or (A3 and A2 and A1 and not(A0) and B3 and not(B2) and B1 and not(B0)) or (A3 and A2 and A1 and not(A0) and B3 and B2 and B1 and B0) or (A3 and A2 and A1 and A0 and B3 and not(B2) and not(B1) and not(B0)) or (A3 and A2 and A1 and A0 and B3 and not(B2) and not(B1) and B0) or (A3 and A2 and A1 and A0 and B3 and not(B2) and B1 and not(B0)) or (A3 and A2 and A1 and A0 and B3 and not(B2) and B1 and B0);
R1 <= (not(A3) and not(A2) and A1 and not(A0) and not(B3) and not(B2) and B1 and B0) or (not(A3) and not(A2) and A1 and not(A0) and not(B3) and B2 and not(B1) and not(B0)) or (not(A3) and not(A2) and A1 and not(A0) and not(B3) and B2 and not(B1) and B0) or (not(A3) and not(A2) and A1 and not(A0) and not(B3) and B2 and B1 and not(B0)) or (not(A3) and not(A2) and A1 and not(A0) and not(B3) and B2 and B1 and B0) or (not(A3) and not(A2) and A1 and not(A0) and B3 and not(B2) and not(B1) and not(B0)) or (not(A3) and not(A2) and A1 and not(A0) and B3 and not(B2) and not(B1) and B0) or (not(A3) and not(A2) and A1 and not(A0) and B3 and not(B2) and B1 and not(B0)) or (not(A3) and not(A2) and A1 and not(A0) and B3 and not(B2) and B1 and B0) or (not(A3) and not(A2) and A1 and not(A0) and B3 and B2 and not(B1) and not(B0)) or (not(A3) and not(A2) and A1 and not(A0) and B3 and B2 and not(B1) and B0) or (not(A3) and not(A2) and A1 and not(A0) and B3 and B2 and B1 and not(B0)) or (not(A3) and not(A2) and A1 and not(A0) and B3 and B2 and B1 and B0) or (not(A3) and not(A2) and A1 and A0 and not(B3) and B2 and not(B1) and not(B0)) or (not(A3) and not(A2) and A1 and A0 and not(B3) and B2 and not(B1) and B0) or (not(A3) and not(A2) and A1 and A0 and not(B3) and B2 and B1 and not(B0)) or (not(A3) and not(A2) and A1 and A0 and not(B3) and B2 and B1 and B0) or (not(A3) and not(A2) and A1 and A0 and B3 and not(B2) and not(B1) and not(B0)) or (not(A3) and not(A2) and A1 and A0 and B3 and not(B2) and not(B1) and B0) or (not(A3) and not(A2) and A1 and A0 and B3 and not(B2) and B1 and not(B0)) or (not(A3) and not(A2) and A1 and A0 and B3 and not(B2) and B1 and B0) or (not(A3) and not(A2) and A1 and A0 and B3 and B2 and not(B1) and not(B0)) or (not(A3) and not(A2) and A1 and A0 and B3 and B2 and not(B1) and B0) or (not(A3) and not(A2) and A1 and A0 and B3 and B2 and B1 and not(B0)) or (not(A3) and not(A2) and A1 and A0 and B3 and B2 and B1 and B0) or (not(A3) and A2 and not(A1) and A0 and not(B3) and not(B2) and B1 and B0) or (not(A3) and A2 and A1 and not(A0) and not(B3) and B2 and not(B1) and not(B0)) or (not(A3) and A2 and A1 and not(A0) and not(B3) and B2 and B1 and B0) or (not(A3) and A2 and A1 and not(A0) and B3 and not(B2) and not(B1) and not(B0)) or (not(A3) and A2 and A1 and not(A0) and B3 and not(B2) and not(B1) and B0) or (not(A3) and A2 and A1 and not(A0) and B3 and not(B2) and B1 and not(B0)) or (not(A3) and A2 and A1 and not(A0) and B3 and not(B2) and B1 and B0) or (not(A3) and A2 and A1 and not(A0) and B3 and B2 and not(B1) and not(B0)) or (not(A3) and A2 and A1 and not(A0) and B3 and B2 and not(B1) and B0) or (not(A3) and A2 and A1 and not(A0) and B3 and B2 and B1 and not(B0)) or (not(A3) and A2 and A1 and not(A0) and B3 and B2 and B1 and B0) or (not(A3) and A2 and A1 and A0 and not(B3) and B2 and not(B1) and not(B0)) or (not(A3) and A2 and A1 and A0 and not(B3) and B2 and not(B1) and B0) or (not(A3) and A2 and A1 and A0 and B3 and not(B2) and not(B1) and not(B0)) or (not(A3) and A2 and A1 and A0 and B3 and not(B2) and not(B1) and B0) or (not(A3) and A2 and A1 and A0 and B3 and not(B2) and B1 and not(B0)) or (not(A3) and A2 and A1 and A0 and B3 and not(B2) and B1 and B0) or (not(A3) and A2 and A1 and A0 and B3 and B2 and not(B1) and not(B0)) or (not(A3) and A2 and A1 and A0 and B3 and B2 and not(B1) and B0) or (not(A3) and A2 and A1 and A0 and B3 and B2 and B1 and not(B0)) or (not(A3) and A2 and A1 and A0 and B3 and B2 and B1 and B0) or (A3 and not(A2) and not(A1) and not(A0) and not(B3) and not(B2) and B1 and B0) or (A3 and not(A2) and not(A1) and not(A0) and not(B3) and B2 and not(B1) and B0) or (A3 and not(A2) and not(A1) and not(A0) and not(B3) and B2 and B1 and not(B0)) or (A3 and not(A2) and not(A1) and A0 and not(B3) and B2 and B1 and not(B0)) or (A3 and not(A2) and not(A1) and A0 and not(B3) and B2 and B1 and B0) or (A3 and not(A2) and A1 and not(A0) and not(B3) and B2 and not(B1) and not(B0)) or (A3 and not(A2) and A1 and not(A0) and not(B3) and B2 and B1 and B0) or (A3 and not(A2) and A1 and not(A0) and B3 and not(B2) and not(B1) and not(B0)) or (A3 and not(A2) and A1 and not(A0) and B3 and not(B2) and B1 and B0) or (A3 and not(A2) and A1 and not(A0) and B3 and B2 and not(B1) and not(B0)) or (A3 and not(A2) and A1 and not(A0) and B3 and B2 and not(B1) and B0) or (A3 and not(A2) and A1 and not(A0) and B3 and B2 and B1 and not(B0)) or (A3 and not(A2) and A1 and not(A0) and B3 and B2 and B1 and B0) or (A3 and not(A2) and A1 and A0 and not(B3) and not(B2) and B1 and B0) or (A3 and not(A2) and A1 and A0 and not(B3) and B2 and not(B1) and not(B0)) or (A3 and not(A2) and A1 and A0 and B3 and not(B2) and not(B1) and not(B0)) or (A3 and not(A2) and A1 and A0 and B3 and not(B2) and not(B1) and B0) or (A3 and not(A2) and A1 and A0 and B3 and B2 and not(B1) and not(B0)) or (A3 and not(A2) and A1 and A0 and B3 and B2 and not(B1) and B0) or (A3 and not(A2) and A1 and A0 and B3 and B2 and B1 and not(B0)) or (A3 and not(A2) and A1 and A0 and B3 and B2 and B1 and B0) or (A3 and A2 and not(A1) and not(A0) and not(B3) and B2 and not(B1) and B0) or (A3 and A2 and not(A1) and not(A0) and B3 and not(B2) and not(B1) and B0) or (A3 and A2 and not(A1) and not(A0) and B3 and not(B2) and B1 and not(B0)) or (A3 and A2 and not(A1) and A0 and not(B3) and B2 and not(B1) and B0) or (A3 and A2 and not(A1) and A0 and not(B3) and B2 and B1 and B0) or (A3 and A2 and not(A1) and A0 and B3 and not(B2) and B1 and not(B0)) or (A3 and A2 and not(A1) and A0 and B3 and not(B2) and B1 and B0) or (A3 and A2 and A1 and not(A0) and not(B3) and not(B2) and B1 and B0) or (A3 and A2 and A1 and not(A0) and not(B3) and B2 and not(B1) and not(B0)) or (A3 and A2 and A1 and not(A0) and not(B3) and B2 and B1 and not(B0)) or (A3 and A2 and A1 and not(A0) and B3 and not(B2) and not(B1) and not(B0)) or (A3 and A2 and A1 and not(A0) and B3 and not(B2) and B1 and B0) or (A3 and A2 and A1 and not(A0) and B3 and B2 and not(B1) and not(B0)) or (A3 and A2 and A1 and not(A0) and B3 and B2 and B1 and B0) or (A3 and A2 and A1 and A0 and not(B3) and B2 and not(B1) and not(B0)) or (A3 and A2 and A1 and A0 and not(B3) and B2 and B1 and not(B0)) or (A3 and A2 and A1 and A0 and B3 and not(B2) and not(B1) and not(B0)) or (A3 and A2 and A1 and A0 and B3 and not(B2) and not(B1) and B0) or (A3 and A2 and A1 and A0 and B3 and B2 and not(B1) and not(B0)) or (A3 and A2 and A1 and A0 and B3 and B2 and not(B1) and B0);
R0 <= (not(A3) and not(A2) and not(A1) and A0 and not(B3) and not(B2) and B1 and not(B0)) or (not(A3) and not(A2) and not(A1) and A0 and not(B3) and not(B2) and B1 and B0) or (not(A3) and not(A2) and not(A1) and A0 and not(B3) and B2 and not(B1) and not(B0)) or (not(A3) and not(A2) and not(A1) and A0 and not(B3) and B2 and not(B1) and B0) or (not(A3) and not(A2) and not(A1) and A0 and not(B3) and B2 and B1 and not(B0)) or (not(A3) and not(A2) and not(A1) and A0 and not(B3) and B2 and B1 and B0) or (not(A3) and not(A2) and not(A1) and A0 and B3 and not(B2) and not(B1) and not(B0)) or (not(A3) and not(A2) and not(A1) and A0 and B3 and not(B2) and not(B1) and B0) or (not(A3) and not(A2) and not(A1) and A0 and B3 and not(B2) and B1 and not(B0)) or (not(A3) and not(A2) and not(A1) and A0 and B3 and not(B2) and B1 and B0) or (not(A3) and not(A2) and not(A1) and A0 and B3 and B2 and not(B1) and not(B0)) or (not(A3) and not(A2) and not(A1) and A0 and B3 and B2 and not(B1) and B0) or (not(A3) and not(A2) and not(A1) and A0 and B3 and B2 and B1 and not(B0)) or (not(A3) and not(A2) and not(A1) and A0 and B3 and B2 and B1 and B0) or (not(A3) and not(A2) and A1 and A0 and not(B3) and not(B2) and B1 and not(B0)) or (not(A3) and not(A2) and A1 and A0 and not(B3) and B2 and not(B1) and not(B0)) or (not(A3) and not(A2) and A1 and A0 and not(B3) and B2 and not(B1) and B0) or (not(A3) and not(A2) and A1 and A0 and not(B3) and B2 and B1 and not(B0)) or (not(A3) and not(A2) and A1 and A0 and not(B3) and B2 and B1 and B0) or (not(A3) and not(A2) and A1 and A0 and B3 and not(B2) and not(B1) and not(B0)) or (not(A3) and not(A2) and A1 and A0 and B3 and not(B2) and not(B1) and B0) or (not(A3) and not(A2) and A1 and A0 and B3 and not(B2) and B1 and not(B0)) or (not(A3) and not(A2) and A1 and A0 and B3 and not(B2) and B1 and B0) or (not(A3) and not(A2) and A1 and A0 and B3 and B2 and not(B1) and not(B0)) or (not(A3) and not(A2) and A1 and A0 and B3 and B2 and not(B1) and B0) or (not(A3) and not(A2) and A1 and A0 and B3 and B2 and B1 and not(B0)) or (not(A3) and not(A2) and A1 and A0 and B3 and B2 and B1 and B0) or (not(A3) and A2 and not(A1) and not(A0) and not(B3) and not(B2) and B1 and B0) or (not(A3) and A2 and not(A1) and A0 and not(B3) and not(B2) and B1 and not(B0)) or (not(A3) and A2 and not(A1) and A0 and not(B3) and B2 and not(B1) and not(B0)) or (not(A3) and A2 and not(A1) and A0 and not(B3) and B2 and B1 and not(B0)) or (not(A3) and A2 and not(A1) and A0 and not(B3) and B2 and B1 and B0) or (not(A3) and A2 and not(A1) and A0 and B3 and not(B2) and not(B1) and not(B0)) or (not(A3) and A2 and not(A1) and A0 and B3 and not(B2) and not(B1) and B0) or (not(A3) and A2 and not(A1) and A0 and B3 and not(B2) and B1 and not(B0)) or (not(A3) and A2 and not(A1) and A0 and B3 and not(B2) and B1 and B0) or (not(A3) and A2 and not(A1) and A0 and B3 and B2 and not(B1) and not(B0)) or (not(A3) and A2 and not(A1) and A0 and B3 and B2 and not(B1) and B0) or (not(A3) and A2 and not(A1) and A0 and B3 and B2 and B1 and not(B0)) or (not(A3) and A2 and not(A1) and A0 and B3 and B2 and B1 and B0) or (not(A3) and A2 and A1 and not(A0) and not(B3) and B2 and not(B1) and B0) or (not(A3) and A2 and A1 and A0 and not(B3) and not(B2) and B1 and not(B0)) or (not(A3) and A2 and A1 and A0 and not(B3) and not(B2) and B1 and B0) or (not(A3) and A2 and A1 and A0 and not(B3) and B2 and not(B1) and not(B0)) or (not(A3) and A2 and A1 and A0 and not(B3) and B2 and B1 and not(B0)) or (not(A3) and A2 and A1 and A0 and B3 and not(B2) and not(B1) and not(B0)) or (not(A3) and A2 and A1 and A0 and B3 and not(B2) and not(B1) and B0) or (not(A3) and A2 and A1 and A0 and B3 and not(B2) and B1 and not(B0)) or (not(A3) and A2 and A1 and A0 and B3 and not(B2) and B1 and B0) or (not(A3) and A2 and A1 and A0 and B3 and B2 and not(B1) and not(B0)) or (not(A3) and A2 and A1 and A0 and B3 and B2 and not(B1) and B0) or (not(A3) and A2 and A1 and A0 and B3 and B2 and B1 and not(B0)) or (not(A3) and A2 and A1 and A0 and B3 and B2 and B1 and B0) or (A3 and not(A2) and not(A1) and not(A0) and not(B3) and B2 and not(B1) and B0) or (A3 and not(A2) and not(A1) and not(A0) and not(B3) and B2 and B1 and B0) or (A3 and not(A2) and not(A1) and A0 and not(B3) and not(B2) and B1 and not(B0)) or (A3 and not(A2) and not(A1) and A0 and not(B3) and B2 and not(B1) and not(B0)) or (A3 and not(A2) and not(A1) and A0 and not(B3) and B2 and B1 and not(B0)) or (A3 and not(A2) and not(A1) and A0 and B3 and not(B2) and not(B1) and not(B0)) or (A3 and not(A2) and not(A1) and A0 and B3 and not(B2) and B1 and not(B0)) or (A3 and not(A2) and not(A1) and A0 and B3 and not(B2) and B1 and B0) or (A3 and not(A2) and not(A1) and A0 and B3 and B2 and not(B1) and not(B0)) or (A3 and not(A2) and not(A1) and A0 and B3 and B2 and not(B1) and B0) or (A3 and not(A2) and not(A1) and A0 and B3 and B2 and B1 and not(B0)) or (A3 and not(A2) and not(A1) and A0 and B3 and B2 and B1 and B0) or (A3 and not(A2) and A1 and not(A0) and not(B3) and not(B2) and B1 and B0) or (A3 and not(A2) and A1 and not(A0) and not(B3) and B2 and B1 and B0) or (A3 and not(A2) and A1 and not(A0) and B3 and not(B2) and not(B1) and B0) or (A3 and not(A2) and A1 and A0 and not(B3) and not(B2) and B1 and not(B0)) or (A3 and not(A2) and A1 and A0 and not(B3) and B2 and not(B1) and not(B0)) or (A3 and not(A2) and A1 and A0 and not(B3) and B2 and not(B1) and B0) or (A3 and not(A2) and A1 and A0 and not(B3) and B2 and B1 and not(B0)) or (A3 and not(A2) and A1 and A0 and B3 and not(B2) and not(B1) and not(B0)) or (A3 and not(A2) and A1 and A0 and B3 and not(B2) and B1 and not(B0)) or (A3 and not(A2) and A1 and A0 and B3 and B2 and not(B1) and not(B0)) or (A3 and not(A2) and A1 and A0 and B3 and B2 and not(B1) and B0) or (A3 and not(A2) and A1 and A0 and B3 and B2 and B1 and not(B0)) or (A3 and not(A2) and A1 and A0 and B3 and B2 and B1 and B0) or (A3 and A2 and not(A1) and not(A0) and not(B3) and B2 and B1 and B0) or (A3 and A2 and not(A1) and not(A0) and B3 and not(B2) and not(B1) and B0) or (A3 and A2 and not(A1) and not(A0) and B3 and not(B2) and B1 and B0) or (A3 and A2 and not(A1) and A0 and not(B3) and not(B2) and B1 and not(B0)) or (A3 and A2 and not(A1) and A0 and not(B3) and not(B2) and B1 and B0) or (A3 and A2 and not(A1) and A0 and not(B3) and B2 and not(B1) and not(B0)) or (A3 and A2 and not(A1) and A0 and not(B3) and B2 and not(B1) and B0) or (A3 and A2 and not(A1) and A0 and not(B3) and B2 and B1 and not(B0)) or (A3 and A2 and not(A1) and A0 and B3 and not(B2) and not(B1) and not(B0)) or (A3 and A2 and not(A1) and A0 and B3 and not(B2) and B1 and not(B0)) or (A3 and A2 and not(A1) and A0 and B3 and B2 and not(B1) and not(B0)) or (A3 and A2 and not(A1) and A0 and B3 and B2 and B1 and not(B0)) or (A3 and A2 and not(A1) and A0 and B3 and B2 and B1 and B0) or (A3 and A2 and A1 and not(A0) and B3 and not(B2) and not(B1) and B0) or (A3 and A2 and A1 and not(A0) and B3 and not(B2) and B1 and B0) or (A3 and A2 and A1 and not(A0) and B3 and B2 and not(B1) and B0) or (A3 and A2 and A1 and A0 and not(B3) and not(B2) and B1 and not(B0)) or (A3 and A2 and A1 and A0 and not(B3) and B2 and not(B1) and not(B0)) or (A3 and A2 and A1 and A0 and not(B3) and B2 and B1 and not(B0)) or (A3 and A2 and A1 and A0 and not(B3) and B2 and B1 and B0) or (A3 and A2 and A1 and A0 and B3 and not(B2) and not(B1) and not(B0)) or (A3 and A2 and A1 and A0 and B3 and not(B2) and B1 and not(B0)) or (A3 and A2 and A1 and A0 and B3 and B2 and not(B1) and not(B0)) or (A3 and A2 and A1 and A0 and B3 and B2 and B1 and not(B0));
end Behavioral;

